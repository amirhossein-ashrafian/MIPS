module AND(
    input a,
    input b,
    output result
);
result = and(result , a, b) ; 
endmodule
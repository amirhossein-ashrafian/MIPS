module MIPS8(
    .input clk ; 
    .input reset ; 
);

endmodule
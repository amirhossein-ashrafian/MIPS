module InstructionMemory (
    input wire clk,                   
    input wire [31:0] PC,       
    output reg [31:0] instruction    
);
    reg [31:0] mem [0:25]; // 26 دستورالعمل

    initial begin

        // برنامه فیبوناچی 

    // دستور lw $0, 0($0)
    mem[0] = 32'b100011_00000_00000_0000000000000000; // opcode:100011 (lw), rs:00000 ($0), rt:00000 ($0), offset:0x0000
    
    // دستور lw $1, 4($0)
    mem[1] = 32'b100011_00000_00001_0000000000000100; // opcode:100011, rs:00000 ($0), rt:00001 ($1), offset:0x0004
    
    // add $2, $0, $1
    mem[2] = 32'b000000_00000_00001_00010_00000_100000; // opcode:000000 (R-type), rs:00000 ($0), rt:00001 ($1), rd:00010 ($2), shamt:00000, funct:100000 (ADD)

    // add $3, $1, $2
    mem[3] = 32'b000000_00001_00010_00011_00000_100000; // rs:00001 ($1), rt:00010 ($2), rd:00011 ($3)

    // add $4, $2, $3
    mem[4] = 32'b000000_00010_00011_00100_00000_100000; // rs:00010 ($2), rt:00011 ($3), rd:00100 ($4)

    // add $5, $3, $4
    mem[5] = 32'b000000_00011_00100_00101_00000_100000; // rs:00011 ($3), rt:00100 ($4), rd:00101 ($5)

    // add $6, $4, $5
    mem[6] = 32'b000000_00100_00101_00110_00000_100000; // rs:00100 ($4), rt:00101 ($5), rd:00110 ($6)

    // add $7, $5, $6
    mem[7] = 32'b000000_00101_00110_00111_00000_100000; // rs:00101 ($5), rt:00110 ($6), rd:00111 ($7)

    // add $8, $6, $7
    mem[8] = 32'b000000_00110_00111_01000_00000_100000; // rs:00110 ($6), rt:00111 ($7), rd:01000 ($8)

    // add $9, $7, $8
    mem[9] = 32'b000000_00111_01000_01001_00000_100000; // rs:00111 ($7), rt:01000 ($8), rd:01001 ($9)

    // add $10, $8, $9
    mem[10] = 32'b000000_01000_01001_01010_00000_100000; // rs:01000 ($8), rt:01001 ($9), rd:01010 ($10)

    // add $11, $9, $10
    mem[11] = 32'b000000_01001_01010_01011_00000_100000; // rs:01001 ($9), rt:01010 ($10), rd:01011 ($11)
    
    // sw $0, 0($0)
    mem[12] = 32'b101011_00000_00000_0000000000000000; // opcode:101011 (sw), rs:00000 ($0), rt:00000 ($0), offset:0x0000

    // sw $1, 4($0)
    mem[13] = 32'b101011_00000_00001_0000000000000100; // rt:00001 ($1), offset:0x0004

    // sw $2, 8($0)
    mem[14] = 32'b101011_00000_00010_0000000000001000; // rt:00010 ($2), offset:0x0008

    // sw $3, 12($0)
    mem[15] = 32'b101011_00000_00011_0000000000001100; // rt:00011 ($3), offset:0x000C

    // sw $4, 16($0)
    mem[16] = 32'b101011_00000_00100_0000000000010000; // rt:00100 ($4), offset:0x0010

    // sw $5, 20($0)
    mem[17] = 32'b101011_00000_00101_0000000000010100; // rt:00101 ($5), offset:0x0014

    // sw $6, 24($0)
    mem[18] = 32'b101011_00000_00110_0000000000011000; // rt:00110 ($6), offset:0x0018

    // sw $7, 28($0)
    mem[19] = 32'b101011_00000_00111_0000000000011100; // rt:00111 ($7), offset:0x001C

    // sw $8, 32($0)
    mem[20] = 32'b101011_00000_01000_0000000000100000; // rt:01000 ($8), offset:0x0020

    // sw $9, 36($0)
    mem[21] = 32'b101011_00000_01001_0000000000100100; // rt:01001 ($9), offset:0x0024

    // sw $10, 40($0)
    mem[22] = 32'b101011_00000_01010_0000000000101000; // rt:01010 ($10), offset:0x0028

    // sw $11, 44($0)
    mem[23] = 32'b101011_00000_01011_0000000000101100; // rt:01011 ($11), offset:0x002C
    end

    always @(posedge clk) begin
        instruction <= mem[PC[31:2]];
    end
endmodule